module reg_write_read();

	test_bench top();
           	reg[31:0] register_tmp;

           	//address
              	parameter TCR_OFFSET   = 12'h00;
              	parameter TDR0_OFFSET  = 12'h04;
              	parameter TDR1_OFFSET  = 12'h08;
              	parameter TCMP0_OFFSET = 12'h0C;
              	parameter TCMP1_OFFSET = 12'h10;
              	parameter TIER_OFFSET  = 12'h14;
              	parameter TISR_OFFSET  = 12'h18;
              	parameter THCSR_OFFSET = 12'h1C;

		initial begin
			#100;				
			$display("\n=======================================TEST WRITE-READ TCR===========================\n");
			top.write(TCR_OFFSET  	, 32'h2222_2222)	;
			top.verify(TCR_OFFSET  	, 32'h0000_0202 )  	;

			$display("\n=================================================END======================================\n");
			
			$display("\n=======================================TEST WRITE-READ TCR===========================\n");
			top.write(TCR_OFFSET  	, 32'h0)	;
			top.verify(TCR_OFFSET  	, 32'h0 )  	;
			$display("\n=================================================END======================================\n");

			$display("\n=======================================TEST WRITE-READ TCR===========================\n");
			top.write(TCR_OFFSET  	, 32'hffff_ffff)	;
			top.verify(TCR_OFFSET  	, 32'h3 )  	;

			$display("\n=================================================END======================================\n");
			
			$display("\n=======================================TEST WRITE-READ TCR===========================\n");
			top.write(TCR_OFFSET  	, 32'h5555_5555)	;
			top.verify(TCR_OFFSET  	, 32'h0000_0501 )  	;
			$display("\n=================================================END======================================\n");

			$display("\n=======================================TEST WRITE-READ TCR===========================\n");
			top.write(TCR_OFFSET  	, 32'hAAAA_AAAA)	;
			top.verify(TCR_OFFSET  	, 32'h0000_0502 )  	;

			$display("\n=================================================END======================================\n");
			
			$display("\n=======================================TEST WRITE-READ TCR===========================\n");
			top.write(TCR_OFFSET  	, 32'h5AA5_A55A)	;
			top.verify(TCR_OFFSET  	, 32'h0000_0502 )  	;
			$display("\n=================================================END======================================\n");

			$display("\n=======================================TEST WRITE-READ TCR===========================\n");
			top.write(TCR_OFFSET  	, 32'h2222_2822)	;
			top.verify(TCR_OFFSET  	, 32'h0000_0802 )  	;

			$display("\n=================================================END======================================\n");
			
			$display("\n=======================================TEST WRITE-READ TCR===========================\n");
			top.write(TCR_OFFSET  	, 32'h2222_2922)	;
			top.verify(TCR_OFFSET  	, 32'h0000_0802 )  	;
			$display("\n=================================================END======================================\n");


			$display("\n=======================================TEST WRITE-READ TCR===========================\n");
			top.write(TCR_OFFSET  	, 32'h2222_2722)	;
			top.verify(TCR_OFFSET  	, 32'h0000_0702 )  	;

			$display("\n=================================================END======================================\n");
			
			$display("\n=======================================TEST WRITE-READ TCR===========================\n");
			top.write(TCR_OFFSET  	, 32'h2222_2622)	;
			top.verify(TCR_OFFSET  	, 32'h0000_0602 )  	;
			$display("\n=================================================END======================================\n");

			$display("\n=======================================TEST WRITE-READ TCR===========================\n");
			top.write(TCR_OFFSET  	, 32'h2222_2422)	;
			top.verify(TCR_OFFSET  	, 32'h0000_0402 )  	;

			$display("\n=================================================END======================================\n");
			
			$display("\n=======================================TEST WRITE-READ TCR===========================\n");
			top.write(TCR_OFFSET  	, 32'h2222_2122)	;
			top.verify(TCR_OFFSET  	, 32'h0000_0102 )  	;
			$display("\n=================================================END======================================\n");






























































			$display("\n=======================================TEST WRITE-READ TDR0===========================\n");
			top.write(TDR0_OFFSET 	, 32'h3333_3333)	;
			top.verify(TDR0_OFFSET 	, 32'h3333_3333)  	;

			$display("\n=================================================END======================================\n");
		
			$display("\n=======================================TEST WRITE-READ TDR0===========================\n");
			top.write(TDR0_OFFSET 	, 32'h1111_1111)	;
			top.verify(TDR0_OFFSET 	, 32'h1111_1111)  	;

			$display("\n=================================================END======================================\n");

			$display("\n=======================================TEST WRITE-READ TDR0===========================\n");
			top.write(TDR0_OFFSET 	, 32'h2222_2222)	;
			top.verify(TDR0_OFFSET 	, 32'h2222_2222)  	;

			$display("\n=================================================END======================================\n");

			$display("\n=======================================TEST WRITE-READ TDR0===========================\n");
			top.write(TDR0_OFFSET 	, 32'hAAAA_AAAA)	;
			top.verify(TDR0_OFFSET 	, 32'hAAAA_AAAA)  	;

			$display("\n=================================================END======================================\n");

			$display("\n=======================================TEST WRITE-READ TDR0===========================\n");
			top.write(TDR0_OFFSET 	, 32'h0)	;
			top.verify(TDR0_OFFSET 	, 32'h0)  	;

			$display("\n=================================================END======================================\n");


			$display("\n=======================================TEST WRITE-READ TDR0===========================\n");
			top.write(TDR0_OFFSET 	, 32'h9999_9999)	;
			top.verify(TDR0_OFFSET 	, 32'h9999_9999)  	;

			$display("\n=================================================END======================================\n");


			$display("\n=======================================TEST WRITE-READ TDR0===========================\n");
			top.write(TDR0_OFFSET 	, 32'h7777_7777)	;
			top.verify(TDR0_OFFSET 	, 32'h7777_7777)  	;

			$display("\n=================================================END======================================\n");


			$display("\n=======================================TEST WRITE-READ TDR1===========================\n");
			top.write(TDR1_OFFSET 	, 32'h4444_4444)	;
			top.verify(TDR1_OFFSET 	, 32'h4444_4444)  	;

			$display("\n=================================================END======================================\n");
			
			$display("\n=======================================TEST WRITE-READ TDR1===========================\n");
			top.write(TDR1_OFFSET 	, 32'h0)	;
			top.verify(TDR1_OFFSET 	, 32'h0)  	;

			$display("\n=================================================END======================================\n");

			$display("\n=======================================TEST WRITE-READ TDR1===========================\n");
			top.write(TDR1_OFFSET 	, 32'h4444_AAAA)	;
			top.verify(TDR1_OFFSET 	, 32'h4444_AAAA)  	;

			$display("\n=================================================END======================================\n");

			$display("\n=======================================TEST WRITE-READ TDR1===========================\n");
			top.write(TDR1_OFFSET 	, 32'h9999_9999)	;
			top.verify(TDR1_OFFSET 	, 32'h9999_9999)  	;

			$display("\n=================================================END======================================\n");


			$display("\n=======================================TEST WRITE-READ TDR1===========================\n");
			top.write(TDR1_OFFSET 	, 32'hCCCC_CCCC)	;
			top.verify(TDR1_OFFSET 	, 32'hCCCC_CCCC)  	;

			$display("\n=================================================END======================================\n");


			$display("\n=======================================TEST WRITE-READ TDR1===========================\n");
			top.write(TDR1_OFFSET 	, 32'h1111_2222)	;
			top.verify(TDR1_OFFSET 	, 32'h1111_2222)  	;

			$display("\n=================================================END======================================\n");


			$display("\n=======================================TEST WRITE-READ TDR1===========================\n");
			top.write(TDR1_OFFSET 	, 32'hABCD_1234)	;
			top.verify(TDR1_OFFSET 	, 32'hABCD_1234)  	;

			$display("\n=================================================END======================================\n");


			$display("\n=======================================TEST WRITE-READ TDR1===========================\n");
			top.write(TDR1_OFFSET 	, 32'hFFFF_FF88)	;
			top.verify(TDR1_OFFSET 	, 32'hFFFF_FF88)  	;

			$display("\n=================================================END======================================\n");


			$display("\n=======================================TEST WRITE-READ TDR1===========================\n");
			top.write(TDR1_OFFSET 	, 32'h1234_5678)	;
			top.verify(TDR1_OFFSET 	, 32'h1234_5678)  	;

			$display("\n=================================================END==================================\n");

			$display("\n=======================================TEST WRITE-READ TCMP0===========================\n");
			top.write(TCMP0_OFFSET	, 32'h5555_5555)	;
			top.verify(TCMP0_OFFSET	, 32'h5555_5555)  	;

			$display("\n=================================================END======================================\n");
		
			$display("\n=======================================TEST WRITE-READ TCMP0===========================\n");
			top.write(TCMP0_OFFSET	, 32'h1234_ABCD)	;
			top.verify(TCMP0_OFFSET	, 32'h1234_ABCD)  	;

			$display("\n=================================================END======================================\n");

			$display("\n=======================================TEST WRITE-READ TCMP0===========================\n");
			top.write(TCMP0_OFFSET	, 32'h5568_5725)	;
			top.verify(TCMP0_OFFSET	, 32'h5568_5725)  	;

			$display("\n=================================================END======================================\n");

			$display("\n=======================================TEST WRITE-READ TCMP0===========================\n");
			top.write(TCMP0_OFFSET	, 32'h0)	;
			top.verify(TCMP0_OFFSET	, 32'h0)  	;

			$display("\n=================================================END======================================\n");


			$display("\n=======================================TEST WRITE-READ TCMP1===========================\n");
			top.write(TCMP1_OFFSET	, 32'h6666_6666)	;
			top.verify(TCMP1_OFFSET	, 32'h6666_6666)  	;

			$display("\n=================================================END======================================\n");

			$display("\n=======================================TEST WRITE-READ TCMP1===========================\n");
			top.write(TCMP1_OFFSET	, 32'h1234_6666)	;
			top.verify(TCMP1_OFFSET	, 32'h1234_6666)  	;

			$display("\n=================================================END======================================\n");

			$display("\n=======================================TEST WRITE-READ TCMP1===========================\n");
			top.write(TCMP1_OFFSET	, 32'hCCAA_6666)	;
			top.verify(TCMP1_OFFSET	, 32'hCCAA_6666)  	;

			$display("\n=================================================END======================================\n");

			$display("\n=======================================TEST WRITE-READ TCMP1===========================\n");
			top.write(TCMP1_OFFSET	, 32'h6677_8866)	;
			top.verify(TCMP1_OFFSET	, 32'h6677_8866)  	;

			$display("\n=================================================END======================================\n");

			$display("\n=======================================TEST WRITE-READ TCMP1===========================\n");
			top.write(TCMP1_OFFSET	, 32'h6326_6596)	;
			top.verify(TCMP1_OFFSET	, 32'h6326_6596)  	;

			$display("\n=================================================END======================================\n");




			$display("\n=======================================TEST WRITE-READ TIER===========================\n");
			top.write(TIER_OFFSET 	, 32'h7777_7777)	;
			top.verify(TIER_OFFSET 	, 32'h1)  	;

			$display("\n=================================================END======================================\n");
		

			$display("\n=======================================TEST WRITE-READ TIER===========================\n");
			top.write(TIER_OFFSET 	, 32'h0)	;
			top.verify(TIER_OFFSET 	, 32'h0)  	;

			$display("\n=================================================END======================================\n");



			$display("\n=======================================TEST WRITE-READ TIER===========================\n");
			top.write(TIER_OFFSET 	, 32'h7777_7773)	;
			top.verify(TIER_OFFSET 	, 32'h1)  	;

			$display("\n=================================================END======================================\n");



			$display("\n=======================================TEST WRITE-READ TIER===========================\n");
			top.write(TIER_OFFSET 	, 32'h7777_777D)	;
			top.verify(TIER_OFFSET 	, 32'h1)  	;

			$display("\n=================================================END======================================\n");





			$display("\n=======================================TEST WRITE-READ TISR===========================\n");
			top.write(TISR_OFFSET 	, 32'h1111_1111)	;
			top.verify(TISR_OFFSET 	, 32'h0)  	;

			$display("\n=================================================END======================================\n");
			

			$display("\n=======================================TEST WRITE-READ TISR===========================\n");
			top.write(TISR_OFFSET 	, 32'hACCC_1110)	;
			top.verify(TISR_OFFSET 	, 32'h0)  	;

			$display("\n=================================================END======================================\n");


			$display("\n=======================================TEST WRITE-READ TISR===========================\n");
			top.write(TISR_OFFSET 	, 32'h11EF_6789)	;
			top.verify(TISR_OFFSET 	, 32'h0)  	;

			$display("\n=================================================END======================================\n");


			$display("\n=======================================TEST WRITE-READ TISR===========================\n");
			top.write(TISR_OFFSET 	, 32'h1111_AAFF)	;
			top.verify(TISR_OFFSET 	, 32'h0)  	;

			$display("\n=================================================END======================================\n");




			$display("\n=======================================TEST WRITE-READ THCSR===========================\n");
			top.write(THCSR_OFFSET	, 32'h8888_8888)	;
			top.verify(THCSR_OFFSET	, 32'h0)  	;

			$display("\n=================================================END======================================\n");
		

			$display("\n=======================================TEST WRITE-READ THCSR===========================\n");
			top.write(THCSR_OFFSET	, 32'h1234_FFF8)	;
			top.verify(THCSR_OFFSET	, 32'h0)  	;

			$display("\n=================================================END======================================\n");


			$display("\n=======================================TEST WRITE-READ THCSR===========================\n");
			top.write(THCSR_OFFSET	, 32'h6969_9696)	;
			top.verify(THCSR_OFFSET	, 32'h0)  	;

			$display("\n=================================================END======================================\n");



			$display("\n=======================================TEST WRITE-READ THCSR===========================\n");
			top.write(THCSR_OFFSET	, 32'hCCDE_8885)	;
			top.verify(THCSR_OFFSET	, 32'h1)  	;

			$display("\n=================================================END======================================\n");


			$display("\n=======================================TEST WRITE-READ THCSR===========================\n");
			top.write(THCSR_OFFSET	, 32'h3223_1293)	;
			top.verify(THCSR_OFFSET	, 32'h1)  	;

			$display("\n=================================================END======================================\n");

		end

endmodule
