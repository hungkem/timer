module check_apb();


endmodule
