module check_onehot();

endmodule
